-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpupkg.all;

entity CtrlROM_ROM is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end CtrlROM_ROM;

architecture arch of CtrlROM_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b0b",
     1 => x"8c0b0b0b",
     2 => x"0b81e004",
     3 => x"0b0b0b0b",
     4 => x"8c04ff0d",
     5 => x"80040400",
     6 => x"00000016",
     7 => x"00000000",
     8 => x"0b0b0bba",
     9 => x"d8080b0b",
    10 => x"0bbadc08",
    11 => x"0b0b0bba",
    12 => x"e0080b0b",
    13 => x"0b0b9808",
    14 => x"2d0b0b0b",
    15 => x"bae00c0b",
    16 => x"0b0bbadc",
    17 => x"0c0b0b0b",
    18 => x"bad80c04",
    19 => x"00000000",
    20 => x"00000000",
    21 => x"00000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"72830609",
    26 => x"81058205",
    27 => x"832b2a83",
    28 => x"ffff0652",
    29 => x"0471fc06",
    30 => x"08728306",
    31 => x"09810583",
    32 => x"05101010",
    33 => x"2a81ff06",
    34 => x"520471fd",
    35 => x"060883ff",
    36 => x"ff738306",
    37 => x"09810582",
    38 => x"05832b2b",
    39 => x"09067383",
    40 => x"ffff0673",
    41 => x"83060981",
    42 => x"05820583",
    43 => x"2b0b2b07",
    44 => x"72fc060c",
    45 => x"51510471",
    46 => x"fc06080b",
    47 => x"0b0bb4dc",
    48 => x"73830610",
    49 => x"10050806",
    50 => x"7381ff06",
    51 => x"73830609",
    52 => x"81058305",
    53 => x"1010102b",
    54 => x"0772fc06",
    55 => x"0c515104",
    56 => x"bad87080",
    57 => x"c594278b",
    58 => x"38807170",
    59 => x"8405530c",
    60 => x"81e2048c",
    61 => x"5188c904",
    62 => x"02fc050d",
    63 => x"f880518f",
    64 => x"0bbae80c",
    65 => x"9f0bbaec",
    66 => x"0ca07170",
    67 => x"81055334",
    68 => x"baec08ff",
    69 => x"05baec0c",
    70 => x"baec0880",
    71 => x"25eb38ba",
    72 => x"e808ff05",
    73 => x"bae80cba",
    74 => x"e8088025",
    75 => x"d738800b",
    76 => x"baec0c80",
    77 => x"0bbae80c",
    78 => x"0284050d",
    79 => x"0402f005",
    80 => x"0df88053",
    81 => x"f8a05483",
    82 => x"bf527370",
    83 => x"81055533",
    84 => x"51707370",
    85 => x"81055534",
    86 => x"ff125271",
    87 => x"8025eb38",
    88 => x"fbc0539f",
    89 => x"52a07370",
    90 => x"81055534",
    91 => x"ff125271",
    92 => x"8025f238",
    93 => x"0290050d",
    94 => x"0402f405",
    95 => x"0d74538e",
    96 => x"0bbae808",
    97 => x"258f3882",
    98 => x"bd2dbae8",
    99 => x"08ff05ba",
   100 => x"e80c82ff",
   101 => x"04bae808",
   102 => x"baec0853",
   103 => x"51728a2e",
   104 => x"098106b7",
   105 => x"38715171",
   106 => x"9f24a038",
   107 => x"bae808a0",
   108 => x"2911f880",
   109 => x"115151a0",
   110 => x"7134baec",
   111 => x"088105ba",
   112 => x"ec0cbaec",
   113 => x"08519f71",
   114 => x"25e23880",
   115 => x"0bbaec0c",
   116 => x"bae80881",
   117 => x"05bae80c",
   118 => x"83ef0470",
   119 => x"a02912f8",
   120 => x"80115151",
   121 => x"727134ba",
   122 => x"ec088105",
   123 => x"baec0cba",
   124 => x"ec08a02e",
   125 => x"0981068e",
   126 => x"38800bba",
   127 => x"ec0cbae8",
   128 => x"088105ba",
   129 => x"e80c028c",
   130 => x"050d0402",
   131 => x"e8050d77",
   132 => x"79565688",
   133 => x"0bfc1677",
   134 => x"712c8f06",
   135 => x"54525480",
   136 => x"53727225",
   137 => x"95387153",
   138 => x"fbe01451",
   139 => x"87713481",
   140 => x"14ff1454",
   141 => x"5472f138",
   142 => x"7153f915",
   143 => x"76712c87",
   144 => x"06535171",
   145 => x"802e8b38",
   146 => x"fbe01451",
   147 => x"71713481",
   148 => x"1454728e",
   149 => x"2495388f",
   150 => x"733153fb",
   151 => x"e01451a0",
   152 => x"71348114",
   153 => x"ff145454",
   154 => x"72f13802",
   155 => x"98050d04",
   156 => x"02ec050d",
   157 => x"800bbaf0",
   158 => x"0cf68c08",
   159 => x"f6900871",
   160 => x"882c5654",
   161 => x"81ff0652",
   162 => x"73722588",
   163 => x"38715482",
   164 => x"0bbaf00c",
   165 => x"72882c73",
   166 => x"81ff0654",
   167 => x"55747325",
   168 => x"8b3872ba",
   169 => x"f0088407",
   170 => x"baf00c55",
   171 => x"73842b86",
   172 => x"a0712583",
   173 => x"7131700b",
   174 => x"0b0bb7b8",
   175 => x"0c81712b",
   176 => x"ff05f688",
   177 => x"0cfdfc13",
   178 => x"ff122c78",
   179 => x"8829ff94",
   180 => x"0570812c",
   181 => x"baf00852",
   182 => x"58525551",
   183 => x"52547680",
   184 => x"2e853870",
   185 => x"81075170",
   186 => x"f6940c71",
   187 => x"098105f6",
   188 => x"800c7209",
   189 => x"8105f684",
   190 => x"0c029405",
   191 => x"0d0402f4",
   192 => x"050d7453",
   193 => x"72708105",
   194 => x"5480f52d",
   195 => x"5271802e",
   196 => x"89387151",
   197 => x"82f92d86",
   198 => x"8404810b",
   199 => x"bad80c02",
   200 => x"8c050d04",
   201 => x"02fc050d",
   202 => x"81808051",
   203 => x"c0115170",
   204 => x"fb380284",
   205 => x"050d0402",
   206 => x"fc050d84",
   207 => x"bf5186a4",
   208 => x"2dff1151",
   209 => x"708025f6",
   210 => x"38028405",
   211 => x"0d0402fc",
   212 => x"050dec51",
   213 => x"83710c86",
   214 => x"a42d8271",
   215 => x"0c028405",
   216 => x"0d0402fc",
   217 => x"050dec51",
   218 => x"8a710c86",
   219 => x"b72d8271",
   220 => x"0c028405",
   221 => x"0d0402fc",
   222 => x"050dec51",
   223 => x"92710c86",
   224 => x"b72d8271",
   225 => x"0c028405",
   226 => x"0d04a00b",
   227 => x"ec0c86b7",
   228 => x"2d0480c0",
   229 => x"0bec0c86",
   230 => x"b72d0402",
   231 => x"dc050d80",
   232 => x"59878a2d",
   233 => x"810bec0c",
   234 => x"7a52baf4",
   235 => x"51ac812d",
   236 => x"bad80879",
   237 => x"2e80ee38",
   238 => x"baf80870",
   239 => x"f80c79ff",
   240 => x"12565955",
   241 => x"73792e8b",
   242 => x"38811874",
   243 => x"812a5558",
   244 => x"73f738f7",
   245 => x"18588159",
   246 => x"80752580",
   247 => x"c8387752",
   248 => x"7351848b",
   249 => x"2dbbcc52",
   250 => x"baf451ae",
   251 => x"c02dbad8",
   252 => x"08802e9a",
   253 => x"38bbcc57",
   254 => x"83fc5676",
   255 => x"70840558",
   256 => x"08e80cfc",
   257 => x"16567580",
   258 => x"25f13888",
   259 => x"9504bad8",
   260 => x"08598480",
   261 => x"55baf451",
   262 => x"ae922dfc",
   263 => x"80158115",
   264 => x"555587d8",
   265 => x"04840bec",
   266 => x"0c78802e",
   267 => x"8d38b7bc",
   268 => x"5190822d",
   269 => x"8df92d88",
   270 => x"c004b8a8",
   271 => x"5190822d",
   272 => x"78bad80c",
   273 => x"02a4050d",
   274 => x"0402f005",
   275 => x"0d840bec",
   276 => x"0c8db02d",
   277 => x"89f72d81",
   278 => x"f82d8352",
   279 => x"8d952d81",
   280 => x"5184f02d",
   281 => x"ff125271",
   282 => x"8025f138",
   283 => x"840bec0c",
   284 => x"b5ec5185",
   285 => x"fe2da380",
   286 => x"2dbad808",
   287 => x"802e80e2",
   288 => x"38879b51",
   289 => x"b4d52db7",
   290 => x"bc519082",
   291 => x"2d8de62d",
   292 => x"8a832d90",
   293 => x"922db7d0",
   294 => x"0b80f52d",
   295 => x"b9940870",
   296 => x"81065455",
   297 => x"5371802e",
   298 => x"85387281",
   299 => x"07537381",
   300 => x"2a708106",
   301 => x"51527180",
   302 => x"2e853872",
   303 => x"82075373",
   304 => x"822a7081",
   305 => x"06515271",
   306 => x"802e8538",
   307 => x"72840753",
   308 => x"72fc0c86",
   309 => x"52bad808",
   310 => x"83388452",
   311 => x"71ec0c89",
   312 => x"9004800b",
   313 => x"bad80c02",
   314 => x"90050d04",
   315 => x"71980c04",
   316 => x"ffb008ba",
   317 => x"d80c0481",
   318 => x"0bffb00c",
   319 => x"04800bff",
   320 => x"b00c0402",
   321 => x"f4050d8b",
   322 => x"8504bad8",
   323 => x"0881f02e",
   324 => x"09810689",
   325 => x"38810bb9",
   326 => x"8c0c8b85",
   327 => x"04bad808",
   328 => x"81e02e09",
   329 => x"81068938",
   330 => x"810bb990",
   331 => x"0c8b8504",
   332 => x"bad80852",
   333 => x"b9900880",
   334 => x"2e8838ba",
   335 => x"d8088180",
   336 => x"05527184",
   337 => x"2c728f06",
   338 => x"5353b98c",
   339 => x"08802e99",
   340 => x"38728429",
   341 => x"b8cc0572",
   342 => x"1381712b",
   343 => x"70097308",
   344 => x"06730c51",
   345 => x"53538afb",
   346 => x"04728429",
   347 => x"b8cc0572",
   348 => x"1383712b",
   349 => x"72080772",
   350 => x"0c535380",
   351 => x"0bb9900c",
   352 => x"800bb98c",
   353 => x"0cbb8051",
   354 => x"8c862dba",
   355 => x"d808ff24",
   356 => x"fef83880",
   357 => x"0bbad80c",
   358 => x"028c050d",
   359 => x"0402f805",
   360 => x"0db8cc52",
   361 => x"8f518072",
   362 => x"70840554",
   363 => x"0cff1151",
   364 => x"708025f2",
   365 => x"38028805",
   366 => x"0d0402f0",
   367 => x"050d7551",
   368 => x"89fd2d70",
   369 => x"822cfc06",
   370 => x"b8cc1172",
   371 => x"109e0671",
   372 => x"0870722a",
   373 => x"70830682",
   374 => x"742b7009",
   375 => x"7406760c",
   376 => x"54515657",
   377 => x"53515389",
   378 => x"f72d71ba",
   379 => x"d80c0290",
   380 => x"050d0402",
   381 => x"fc050d72",
   382 => x"5180710c",
   383 => x"800b8412",
   384 => x"0c028405",
   385 => x"0d0402f0",
   386 => x"050d7570",
   387 => x"08841208",
   388 => x"535353ff",
   389 => x"5471712e",
   390 => x"a83889fd",
   391 => x"2d841308",
   392 => x"70842914",
   393 => x"88117008",
   394 => x"7081ff06",
   395 => x"84180881",
   396 => x"11870684",
   397 => x"1a0c5351",
   398 => x"55515151",
   399 => x"89f72d71",
   400 => x"5473bad8",
   401 => x"0c029005",
   402 => x"0d0402f4",
   403 => x"050d89fd",
   404 => x"2de00870",
   405 => x"8b2a7081",
   406 => x"06515253",
   407 => x"70802e9d",
   408 => x"38bb8008",
   409 => x"708429bb",
   410 => x"88057481",
   411 => x"ff06710c",
   412 => x"5151bb80",
   413 => x"08811187",
   414 => x"06bb800c",
   415 => x"51728c2c",
   416 => x"bf06bba8",
   417 => x"0c800bbb",
   418 => x"ac0c89f0",
   419 => x"2d89f72d",
   420 => x"028c050d",
   421 => x"0402fc05",
   422 => x"0d89fd2d",
   423 => x"810bbbac",
   424 => x"0c89f72d",
   425 => x"bbac0851",
   426 => x"70fa3802",
   427 => x"84050d04",
   428 => x"02fc050d",
   429 => x"bb80518b",
   430 => x"f32d8b9d",
   431 => x"2d8cca51",
   432 => x"89ec2d02",
   433 => x"84050d04",
   434 => x"02fc050d",
   435 => x"8fcf5186",
   436 => x"a42dff11",
   437 => x"51708025",
   438 => x"f6380284",
   439 => x"050d04bb",
   440 => x"b808bad8",
   441 => x"0c0402fc",
   442 => x"050d810b",
   443 => x"b9980c81",
   444 => x"5184f02d",
   445 => x"0284050d",
   446 => x"0402f805",
   447 => x"0d8e8304",
   448 => x"8a832d80",
   449 => x"f6518bba",
   450 => x"2dbad808",
   451 => x"f33880da",
   452 => x"518bba2d",
   453 => x"bad808e8",
   454 => x"38bba808",
   455 => x"80c00652",
   456 => x"718024dc",
   457 => x"38bad808",
   458 => x"b9980cba",
   459 => x"d8085184",
   460 => x"f02d0288",
   461 => x"050d0402",
   462 => x"ec050d76",
   463 => x"54805287",
   464 => x"0b881580",
   465 => x"f52d5653",
   466 => x"74722483",
   467 => x"38a05372",
   468 => x"5182f92d",
   469 => x"81128b15",
   470 => x"80f52d54",
   471 => x"52727225",
   472 => x"de380294",
   473 => x"050d0402",
   474 => x"f0050dbb",
   475 => x"b8085481",
   476 => x"f82d800b",
   477 => x"bbbc0c73",
   478 => x"08802e81",
   479 => x"8038820b",
   480 => x"baec0cbb",
   481 => x"bc088f06",
   482 => x"bae80c73",
   483 => x"08527183",
   484 => x"2e963871",
   485 => x"83268938",
   486 => x"71812eaf",
   487 => x"388fe804",
   488 => x"71852e9f",
   489 => x"388fe804",
   490 => x"881480f5",
   491 => x"2d841508",
   492 => x"b6845354",
   493 => x"5285fe2d",
   494 => x"71842913",
   495 => x"70085252",
   496 => x"8fec0473",
   497 => x"518eb72d",
   498 => x"8fe804b9",
   499 => x"94088815",
   500 => x"082c7081",
   501 => x"06515271",
   502 => x"802e8738",
   503 => x"b688518f",
   504 => x"e504b68c",
   505 => x"5185fe2d",
   506 => x"84140851",
   507 => x"85fe2dbb",
   508 => x"bc088105",
   509 => x"bbbc0c8c",
   510 => x"14548ef7",
   511 => x"04029005",
   512 => x"0d0471bb",
   513 => x"b80c8ee7",
   514 => x"2dbbbc08",
   515 => x"ff05bbc0",
   516 => x"0c0402e8",
   517 => x"050dbbb8",
   518 => x"08bbc408",
   519 => x"575580f6",
   520 => x"518bba2d",
   521 => x"bad80881",
   522 => x"2a708106",
   523 => x"51527193",
   524 => x"38bba808",
   525 => x"80c00652",
   526 => x"8072259f",
   527 => x"3890c304",
   528 => x"8a832d80",
   529 => x"f6518bba",
   530 => x"2dbad808",
   531 => x"f338b998",
   532 => x"08813270",
   533 => x"b9980c51",
   534 => x"84f02dbb",
   535 => x"a808a006",
   536 => x"52807225",
   537 => x"96388dc8",
   538 => x"2d8a832d",
   539 => x"b9980881",
   540 => x"3270b998",
   541 => x"0c705252",
   542 => x"84f02d80",
   543 => x"0bbbb00c",
   544 => x"800bbbb4",
   545 => x"0cb99808",
   546 => x"83b93880",
   547 => x"da518bba",
   548 => x"2dbad808",
   549 => x"802e8a38",
   550 => x"bbb00881",
   551 => x"8007bbb0",
   552 => x"0c80d951",
   553 => x"8bba2dba",
   554 => x"d808802e",
   555 => x"8a38bbb0",
   556 => x"0880c007",
   557 => x"bbb00c81",
   558 => x"94518bba",
   559 => x"2dbad808",
   560 => x"802e8938",
   561 => x"bbb00890",
   562 => x"07bbb00c",
   563 => x"8191518b",
   564 => x"ba2dbad8",
   565 => x"08802e89",
   566 => x"38bbb008",
   567 => x"a007bbb0",
   568 => x"0c81f551",
   569 => x"8bba2dba",
   570 => x"d808802e",
   571 => x"8938bbb0",
   572 => x"088107bb",
   573 => x"b00c81f2",
   574 => x"518bba2d",
   575 => x"bad80880",
   576 => x"2e8938bb",
   577 => x"b0088207",
   578 => x"bbb00c81",
   579 => x"eb518bba",
   580 => x"2dbad808",
   581 => x"802e8938",
   582 => x"bbb00884",
   583 => x"07bbb00c",
   584 => x"81f4518b",
   585 => x"ba2dbad8",
   586 => x"08802e89",
   587 => x"38bbb008",
   588 => x"8807bbb0",
   589 => x"0c80d851",
   590 => x"8bba2dba",
   591 => x"d808802e",
   592 => x"8a38bbb4",
   593 => x"08818007",
   594 => x"bbb40c92",
   595 => x"518bba2d",
   596 => x"bad80880",
   597 => x"2e8a38bb",
   598 => x"b40880c0",
   599 => x"07bbb40c",
   600 => x"94518bba",
   601 => x"2dbad808",
   602 => x"802e8938",
   603 => x"bbb40890",
   604 => x"07bbb40c",
   605 => x"91518bba",
   606 => x"2dbad808",
   607 => x"802e8938",
   608 => x"bbb408a0",
   609 => x"07bbb40c",
   610 => x"9d518bba",
   611 => x"2dbad808",
   612 => x"802e8938",
   613 => x"bbb40881",
   614 => x"07bbb40c",
   615 => x"9b518bba",
   616 => x"2dbad808",
   617 => x"802e8938",
   618 => x"bbb40882",
   619 => x"07bbb40c",
   620 => x"9c518bba",
   621 => x"2dbad808",
   622 => x"802e8938",
   623 => x"bbb40884",
   624 => x"07bbb40c",
   625 => x"a3518bba",
   626 => x"2dbad808",
   627 => x"802e8938",
   628 => x"bbb40888",
   629 => x"07bbb40c",
   630 => x"96518bba",
   631 => x"2dbad808",
   632 => x"802e8438",
   633 => x"86f62d9e",
   634 => x"518bba2d",
   635 => x"bad80880",
   636 => x"2e843886",
   637 => x"e22d9451",
   638 => x"8bba2dba",
   639 => x"d8088e38",
   640 => x"8194518b",
   641 => x"ba2dbad8",
   642 => x"08802ea8",
   643 => x"3891518b",
   644 => x"ba2dbad8",
   645 => x"088e3881",
   646 => x"91518bba",
   647 => x"2dbad808",
   648 => x"802e9138",
   649 => x"80e6518b",
   650 => x"ba2dbad8",
   651 => x"08802e84",
   652 => x"3887922d",
   653 => x"81fd518b",
   654 => x"ba2d81fa",
   655 => x"518bba2d",
   656 => x"9af70494",
   657 => x"518bba2d",
   658 => x"bad8088e",
   659 => x"38819451",
   660 => x"8bba2dba",
   661 => x"d808802e",
   662 => x"a8389151",
   663 => x"8bba2dba",
   664 => x"d8088e38",
   665 => x"8191518b",
   666 => x"ba2dbad8",
   667 => x"08802e91",
   668 => x"3880e651",
   669 => x"8bba2dba",
   670 => x"d808802e",
   671 => x"84388792",
   672 => x"2d81f551",
   673 => x"8bba2dba",
   674 => x"d808812a",
   675 => x"70810651",
   676 => x"52718c38",
   677 => x"bba80890",
   678 => x"06528072",
   679 => x"25bd38bb",
   680 => x"a8089006",
   681 => x"52807225",
   682 => x"84388dc8",
   683 => x"2dbbc008",
   684 => x"5271802e",
   685 => x"8938ff12",
   686 => x"bbc00c95",
   687 => x"db04bbbc",
   688 => x"0810bbbc",
   689 => x"08057084",
   690 => x"29165152",
   691 => x"88120880",
   692 => x"2e8938ff",
   693 => x"51881208",
   694 => x"52712d81",
   695 => x"f2518bba",
   696 => x"2dbad808",
   697 => x"812a7081",
   698 => x"06515271",
   699 => x"8c38bba8",
   700 => x"08880652",
   701 => x"807225bf",
   702 => x"38bba808",
   703 => x"88065280",
   704 => x"72258438",
   705 => x"8dc82dbb",
   706 => x"bc08ff11",
   707 => x"bbc00856",
   708 => x"53537372",
   709 => x"25893881",
   710 => x"14bbc00c",
   711 => x"96b70472",
   712 => x"10137084",
   713 => x"29165152",
   714 => x"88120880",
   715 => x"2e8938fe",
   716 => x"51881208",
   717 => x"52712d81",
   718 => x"fd518bba",
   719 => x"2dbad808",
   720 => x"812a7081",
   721 => x"06515271",
   722 => x"802ead38",
   723 => x"bbc00880",
   724 => x"2e893880",
   725 => x"0bbbc00c",
   726 => x"96f804bb",
   727 => x"bc0810bb",
   728 => x"bc080570",
   729 => x"84291651",
   730 => x"52881208",
   731 => x"802e8938",
   732 => x"fd518812",
   733 => x"0852712d",
   734 => x"81fa518b",
   735 => x"ba2dbad8",
   736 => x"08812a70",
   737 => x"81065152",
   738 => x"71802eae",
   739 => x"38bbbc08",
   740 => x"ff115452",
   741 => x"bbc00873",
   742 => x"25883872",
   743 => x"bbc00c97",
   744 => x"ba047110",
   745 => x"12708429",
   746 => x"16515288",
   747 => x"1208802e",
   748 => x"8938fc51",
   749 => x"88120852",
   750 => x"712dbbc0",
   751 => x"08705354",
   752 => x"73802e8a",
   753 => x"388c15ff",
   754 => x"15555597",
   755 => x"c004820b",
   756 => x"baec0c71",
   757 => x"8f06bae8",
   758 => x"0c81eb51",
   759 => x"8bba2dba",
   760 => x"d808812a",
   761 => x"70810651",
   762 => x"5271802e",
   763 => x"ad387408",
   764 => x"852e0981",
   765 => x"06a43888",
   766 => x"1580f52d",
   767 => x"ff055271",
   768 => x"881681b7",
   769 => x"2d71982b",
   770 => x"52718025",
   771 => x"8838800b",
   772 => x"881681b7",
   773 => x"2d74518e",
   774 => x"b72d81f4",
   775 => x"518bba2d",
   776 => x"bad80881",
   777 => x"2a708106",
   778 => x"51527180",
   779 => x"2eb33874",
   780 => x"08852e09",
   781 => x"8106aa38",
   782 => x"881580f5",
   783 => x"2d810552",
   784 => x"71881681",
   785 => x"b72d7181",
   786 => x"ff068b16",
   787 => x"80f52d54",
   788 => x"52727227",
   789 => x"87387288",
   790 => x"1681b72d",
   791 => x"74518eb7",
   792 => x"2d80da51",
   793 => x"8bba2dba",
   794 => x"d808812a",
   795 => x"70810651",
   796 => x"52718d38",
   797 => x"bba80881",
   798 => x"06528072",
   799 => x"2581b438",
   800 => x"bbb808bb",
   801 => x"a8088106",
   802 => x"53538072",
   803 => x"2584388d",
   804 => x"c82dbbc0",
   805 => x"08547380",
   806 => x"2e8a388c",
   807 => x"13ff1555",
   808 => x"53999604",
   809 => x"72085271",
   810 => x"822ea638",
   811 => x"71822689",
   812 => x"3871812e",
   813 => x"a9389ab3",
   814 => x"0471832e",
   815 => x"b1387184",
   816 => x"2e098106",
   817 => x"80ed3888",
   818 => x"13085190",
   819 => x"822d9ab3",
   820 => x"04bbc008",
   821 => x"51881308",
   822 => x"52712d9a",
   823 => x"b304810b",
   824 => x"8814082b",
   825 => x"b9940832",
   826 => x"b9940c9a",
   827 => x"89048813",
   828 => x"80f52d81",
   829 => x"058b1480",
   830 => x"f52d5354",
   831 => x"71742483",
   832 => x"38805473",
   833 => x"881481b7",
   834 => x"2d8ee72d",
   835 => x"9ab30475",
   836 => x"08802ea2",
   837 => x"38750851",
   838 => x"8bba2dba",
   839 => x"d8088106",
   840 => x"5271802e",
   841 => x"8b38bbc0",
   842 => x"08518416",
   843 => x"0852712d",
   844 => x"88165675",
   845 => x"da388054",
   846 => x"800bbaec",
   847 => x"0c738f06",
   848 => x"bae80ca0",
   849 => x"5273bbc0",
   850 => x"082e0981",
   851 => x"069838bb",
   852 => x"bc08ff05",
   853 => x"74327009",
   854 => x"81057072",
   855 => x"079f2a91",
   856 => x"71315151",
   857 => x"53537151",
   858 => x"82f92d81",
   859 => x"14548e74",
   860 => x"25c638b9",
   861 => x"98085271",
   862 => x"bad80c02",
   863 => x"98050d04",
   864 => x"02f4050d",
   865 => x"d45281ff",
   866 => x"720c7108",
   867 => x"5381ff72",
   868 => x"0c72882b",
   869 => x"83fe8006",
   870 => x"72087081",
   871 => x"ff065152",
   872 => x"5381ff72",
   873 => x"0c727107",
   874 => x"882b7208",
   875 => x"7081ff06",
   876 => x"51525381",
   877 => x"ff720c72",
   878 => x"7107882b",
   879 => x"72087081",
   880 => x"ff067207",
   881 => x"bad80c52",
   882 => x"53028c05",
   883 => x"0d0402f4",
   884 => x"050d7476",
   885 => x"7181ff06",
   886 => x"d40c5353",
   887 => x"bbc80885",
   888 => x"3871892b",
   889 => x"5271982a",
   890 => x"d40c7190",
   891 => x"2a7081ff",
   892 => x"06d40c51",
   893 => x"71882a70",
   894 => x"81ff06d4",
   895 => x"0c517181",
   896 => x"ff06d40c",
   897 => x"72902a70",
   898 => x"81ff06d4",
   899 => x"0c51d408",
   900 => x"7081ff06",
   901 => x"515182b8",
   902 => x"bf527081",
   903 => x"ff2e0981",
   904 => x"06943881",
   905 => x"ff0bd40c",
   906 => x"d4087081",
   907 => x"ff06ff14",
   908 => x"54515171",
   909 => x"e53870ba",
   910 => x"d80c028c",
   911 => x"050d0402",
   912 => x"fc050d81",
   913 => x"c75181ff",
   914 => x"0bd40cff",
   915 => x"11517080",
   916 => x"25f43802",
   917 => x"84050d04",
   918 => x"02f4050d",
   919 => x"81ff0bd4",
   920 => x"0c935380",
   921 => x"5287fc80",
   922 => x"c1519bce",
   923 => x"2dbad808",
   924 => x"8b3881ff",
   925 => x"0bd40c81",
   926 => x"539d8504",
   927 => x"9cbf2dff",
   928 => x"135372df",
   929 => x"3872bad8",
   930 => x"0c028c05",
   931 => x"0d0402ec",
   932 => x"050d810b",
   933 => x"bbc80c84",
   934 => x"54d00870",
   935 => x"8f2a7081",
   936 => x"06515153",
   937 => x"72f33872",
   938 => x"d00c9cbf",
   939 => x"2db69051",
   940 => x"85fe2dd0",
   941 => x"08708f2a",
   942 => x"70810651",
   943 => x"515372f3",
   944 => x"38810bd0",
   945 => x"0cb15380",
   946 => x"5284d480",
   947 => x"c0519bce",
   948 => x"2dbad808",
   949 => x"812e9338",
   950 => x"72822ebd",
   951 => x"38ff1353",
   952 => x"72e538ff",
   953 => x"145473ff",
   954 => x"b0389cbf",
   955 => x"2d83aa52",
   956 => x"849c80c8",
   957 => x"519bce2d",
   958 => x"bad80881",
   959 => x"2e098106",
   960 => x"92389b80",
   961 => x"2dbad808",
   962 => x"83ffff06",
   963 => x"537283aa",
   964 => x"2e9d389c",
   965 => x"d82d9eaa",
   966 => x"04b69c51",
   967 => x"85fe2d80",
   968 => x"539ff804",
   969 => x"b6b45185",
   970 => x"fe2d8054",
   971 => x"9fca0481",
   972 => x"ff0bd40c",
   973 => x"b1549cbf",
   974 => x"2d8fcf53",
   975 => x"805287fc",
   976 => x"80f7519b",
   977 => x"ce2dbad8",
   978 => x"0855bad8",
   979 => x"08812e09",
   980 => x"81069b38",
   981 => x"81ff0bd4",
   982 => x"0c820a52",
   983 => x"849c80e9",
   984 => x"519bce2d",
   985 => x"bad80880",
   986 => x"2e8d389c",
   987 => x"bf2dff13",
   988 => x"5372c938",
   989 => x"9fbd0481",
   990 => x"ff0bd40c",
   991 => x"bad80852",
   992 => x"87fc80fa",
   993 => x"519bce2d",
   994 => x"bad808b1",
   995 => x"3881ff0b",
   996 => x"d40cd408",
   997 => x"5381ff0b",
   998 => x"d40c81ff",
   999 => x"0bd40c81",
  1000 => x"ff0bd40c",
  1001 => x"81ff0bd4",
  1002 => x"0c72862a",
  1003 => x"70810676",
  1004 => x"56515372",
  1005 => x"9538bad8",
  1006 => x"08549fca",
  1007 => x"0473822e",
  1008 => x"fee238ff",
  1009 => x"145473fe",
  1010 => x"ed3873bb",
  1011 => x"c80c738b",
  1012 => x"38815287",
  1013 => x"fc80d051",
  1014 => x"9bce2d81",
  1015 => x"ff0bd40c",
  1016 => x"d008708f",
  1017 => x"2a708106",
  1018 => x"51515372",
  1019 => x"f33872d0",
  1020 => x"0c81ff0b",
  1021 => x"d40c8153",
  1022 => x"72bad80c",
  1023 => x"0294050d",
  1024 => x"0402e805",
  1025 => x"0d785580",
  1026 => x"5681ff0b",
  1027 => x"d40cd008",
  1028 => x"708f2a70",
  1029 => x"81065151",
  1030 => x"5372f338",
  1031 => x"82810bd0",
  1032 => x"0c81ff0b",
  1033 => x"d40c7752",
  1034 => x"87fc80d1",
  1035 => x"519bce2d",
  1036 => x"80dbc6df",
  1037 => x"54bad808",
  1038 => x"802e8a38",
  1039 => x"b6d45185",
  1040 => x"fe2da198",
  1041 => x"0481ff0b",
  1042 => x"d40cd408",
  1043 => x"7081ff06",
  1044 => x"51537281",
  1045 => x"fe2e0981",
  1046 => x"069d3880",
  1047 => x"ff539b80",
  1048 => x"2dbad808",
  1049 => x"75708405",
  1050 => x"570cff13",
  1051 => x"53728025",
  1052 => x"ed388156",
  1053 => x"a0fd04ff",
  1054 => x"145473c9",
  1055 => x"3881ff0b",
  1056 => x"d40c81ff",
  1057 => x"0bd40cd0",
  1058 => x"08708f2a",
  1059 => x"70810651",
  1060 => x"515372f3",
  1061 => x"3872d00c",
  1062 => x"75bad80c",
  1063 => x"0298050d",
  1064 => x"0402e805",
  1065 => x"0d77797b",
  1066 => x"58555580",
  1067 => x"53727625",
  1068 => x"a3387470",
  1069 => x"81055680",
  1070 => x"f52d7470",
  1071 => x"81055680",
  1072 => x"f52d5252",
  1073 => x"71712e86",
  1074 => x"388151a1",
  1075 => x"d6048113",
  1076 => x"53a1ad04",
  1077 => x"805170ba",
  1078 => x"d80c0298",
  1079 => x"050d0402",
  1080 => x"ec050d76",
  1081 => x"5574802e",
  1082 => x"be389a15",
  1083 => x"80e02d51",
  1084 => x"af992dba",
  1085 => x"d808bad8",
  1086 => x"0880c1fc",
  1087 => x"0cbad808",
  1088 => x"545480c1",
  1089 => x"d808802e",
  1090 => x"99389415",
  1091 => x"80e02d51",
  1092 => x"af992dba",
  1093 => x"d808902b",
  1094 => x"83fff00a",
  1095 => x"06707507",
  1096 => x"51537280",
  1097 => x"c1fc0c80",
  1098 => x"c1fc0853",
  1099 => x"72802e9d",
  1100 => x"3880c1d0",
  1101 => x"08fe1471",
  1102 => x"2980c1e4",
  1103 => x"080580c2",
  1104 => x"800c7084",
  1105 => x"2b80c1dc",
  1106 => x"0c54a2fb",
  1107 => x"0480c1e8",
  1108 => x"0880c1fc",
  1109 => x"0c80c1ec",
  1110 => x"0880c280",
  1111 => x"0c80c1d8",
  1112 => x"08802e8b",
  1113 => x"3880c1d0",
  1114 => x"08842b53",
  1115 => x"a2f60480",
  1116 => x"c1f00884",
  1117 => x"2b537280",
  1118 => x"c1dc0c02",
  1119 => x"94050d04",
  1120 => x"02d8050d",
  1121 => x"800b80c1",
  1122 => x"d80c8454",
  1123 => x"9d8e2dba",
  1124 => x"d808802e",
  1125 => x"9538bbcc",
  1126 => x"528051a0",
  1127 => x"812dbad8",
  1128 => x"08802e86",
  1129 => x"38fe54a3",
  1130 => x"b204ff14",
  1131 => x"54738024",
  1132 => x"db38738c",
  1133 => x"38b6e451",
  1134 => x"85fe2d73",
  1135 => x"55a8d404",
  1136 => x"8056810b",
  1137 => x"80c2840c",
  1138 => x"8853b6f8",
  1139 => x"52bc8251",
  1140 => x"a1a12dba",
  1141 => x"d808762e",
  1142 => x"09810688",
  1143 => x"38bad808",
  1144 => x"80c2840c",
  1145 => x"8853b784",
  1146 => x"52bc9e51",
  1147 => x"a1a12dba",
  1148 => x"d8088838",
  1149 => x"bad80880",
  1150 => x"c2840c80",
  1151 => x"c2840880",
  1152 => x"2e80f638",
  1153 => x"bf920b80",
  1154 => x"f52dbf93",
  1155 => x"0b80f52d",
  1156 => x"71982b71",
  1157 => x"902b07bf",
  1158 => x"940b80f5",
  1159 => x"2d70882b",
  1160 => x"7207bf95",
  1161 => x"0b80f52d",
  1162 => x"7107bfca",
  1163 => x"0b80f52d",
  1164 => x"bfcb0b80",
  1165 => x"f52d7188",
  1166 => x"2b07535f",
  1167 => x"54525a56",
  1168 => x"57557381",
  1169 => x"abaa2e09",
  1170 => x"81068d38",
  1171 => x"7551aee9",
  1172 => x"2dbad808",
  1173 => x"56a4e504",
  1174 => x"7382d4d5",
  1175 => x"2e8738b7",
  1176 => x"9051a5a7",
  1177 => x"04bbcc52",
  1178 => x"7551a081",
  1179 => x"2dbad808",
  1180 => x"55bad808",
  1181 => x"802e83dc",
  1182 => x"388853b7",
  1183 => x"8452bc9e",
  1184 => x"51a1a12d",
  1185 => x"bad8088a",
  1186 => x"38810b80",
  1187 => x"c1d80ca5",
  1188 => x"ad048853",
  1189 => x"b6f852bc",
  1190 => x"8251a1a1",
  1191 => x"2dbad808",
  1192 => x"802e8a38",
  1193 => x"b7a45185",
  1194 => x"fe2da687",
  1195 => x"04bfca0b",
  1196 => x"80f52d54",
  1197 => x"7380d52e",
  1198 => x"09810680",
  1199 => x"ca38bfcb",
  1200 => x"0b80f52d",
  1201 => x"547381aa",
  1202 => x"2e098106",
  1203 => x"ba38800b",
  1204 => x"bbcc0b80",
  1205 => x"f52d5654",
  1206 => x"7481e92e",
  1207 => x"83388154",
  1208 => x"7481eb2e",
  1209 => x"8c388055",
  1210 => x"73752e09",
  1211 => x"810682e4",
  1212 => x"38bbd70b",
  1213 => x"80f52d55",
  1214 => x"748d38bb",
  1215 => x"d80b80f5",
  1216 => x"2d547382",
  1217 => x"2e863880",
  1218 => x"55a8d404",
  1219 => x"bbd90b80",
  1220 => x"f52d7080",
  1221 => x"c1d00cff",
  1222 => x"0580c1d4",
  1223 => x"0cbbda0b",
  1224 => x"80f52dbb",
  1225 => x"db0b80f5",
  1226 => x"2d587605",
  1227 => x"77828029",
  1228 => x"057080c1",
  1229 => x"e00cbbdc",
  1230 => x"0b80f52d",
  1231 => x"7080c1f4",
  1232 => x"0c80c1d8",
  1233 => x"08595758",
  1234 => x"76802e81",
  1235 => x"ac388853",
  1236 => x"b78452bc",
  1237 => x"9e51a1a1",
  1238 => x"2dbad808",
  1239 => x"81f63880",
  1240 => x"c1d00870",
  1241 => x"842b80c1",
  1242 => x"dc0c7080",
  1243 => x"c1f00cbb",
  1244 => x"f10b80f5",
  1245 => x"2dbbf00b",
  1246 => x"80f52d71",
  1247 => x"82802905",
  1248 => x"bbf20b80",
  1249 => x"f52d7084",
  1250 => x"80802912",
  1251 => x"bbf30b80",
  1252 => x"f52d7081",
  1253 => x"800a2912",
  1254 => x"7080c1f8",
  1255 => x"0c80c1f4",
  1256 => x"08712980",
  1257 => x"c1e00805",
  1258 => x"7080c1e4",
  1259 => x"0cbbf90b",
  1260 => x"80f52dbb",
  1261 => x"f80b80f5",
  1262 => x"2d718280",
  1263 => x"2905bbfa",
  1264 => x"0b80f52d",
  1265 => x"70848080",
  1266 => x"2912bbfb",
  1267 => x"0b80f52d",
  1268 => x"70982b81",
  1269 => x"f00a0672",
  1270 => x"057080c1",
  1271 => x"e80cfe11",
  1272 => x"7e297705",
  1273 => x"80c1ec0c",
  1274 => x"52595243",
  1275 => x"545e5152",
  1276 => x"59525d57",
  1277 => x"5957a8cd",
  1278 => x"04bbde0b",
  1279 => x"80f52dbb",
  1280 => x"dd0b80f5",
  1281 => x"2d718280",
  1282 => x"29057080",
  1283 => x"c1dc0c70",
  1284 => x"a02983ff",
  1285 => x"0570892a",
  1286 => x"7080c1f0",
  1287 => x"0cbbe30b",
  1288 => x"80f52dbb",
  1289 => x"e20b80f5",
  1290 => x"2d718280",
  1291 => x"29057080",
  1292 => x"c1f80c7b",
  1293 => x"71291e70",
  1294 => x"80c1ec0c",
  1295 => x"7d80c1e8",
  1296 => x"0c730580",
  1297 => x"c1e40c55",
  1298 => x"5e515155",
  1299 => x"558051a1",
  1300 => x"df2d8155",
  1301 => x"74bad80c",
  1302 => x"02a8050d",
  1303 => x"0402ec05",
  1304 => x"0d767087",
  1305 => x"2c7180ff",
  1306 => x"06555654",
  1307 => x"80c1d808",
  1308 => x"8a387388",
  1309 => x"2c7481ff",
  1310 => x"065455bb",
  1311 => x"cc5280c1",
  1312 => x"e0081551",
  1313 => x"a0812dba",
  1314 => x"d80854ba",
  1315 => x"d808802e",
  1316 => x"b43880c1",
  1317 => x"d808802e",
  1318 => x"98387284",
  1319 => x"29bbcc05",
  1320 => x"70085253",
  1321 => x"aee92dba",
  1322 => x"d808f00a",
  1323 => x"0653a9c3",
  1324 => x"047210bb",
  1325 => x"cc057080",
  1326 => x"e02d5253",
  1327 => x"af992dba",
  1328 => x"d8085372",
  1329 => x"5473bad8",
  1330 => x"0c029405",
  1331 => x"0d0402e0",
  1332 => x"050d7970",
  1333 => x"842c80c2",
  1334 => x"80080571",
  1335 => x"8f065255",
  1336 => x"53728938",
  1337 => x"bbcc5273",
  1338 => x"51a0812d",
  1339 => x"72a029bb",
  1340 => x"cc055480",
  1341 => x"7480f52d",
  1342 => x"56537473",
  1343 => x"2e833881",
  1344 => x"537481e5",
  1345 => x"2e81ef38",
  1346 => x"81707406",
  1347 => x"54587280",
  1348 => x"2e81e338",
  1349 => x"8b1480f5",
  1350 => x"2d70832a",
  1351 => x"79065856",
  1352 => x"769838b9",
  1353 => x"9c085372",
  1354 => x"883872bf",
  1355 => x"cc0b81b7",
  1356 => x"2d76b99c",
  1357 => x"0c7353ab",
  1358 => x"f804758f",
  1359 => x"2e098106",
  1360 => x"81b43874",
  1361 => x"9f068d29",
  1362 => x"bfbf1151",
  1363 => x"53811480",
  1364 => x"f52d7370",
  1365 => x"81055581",
  1366 => x"b72d8314",
  1367 => x"80f52d73",
  1368 => x"70810555",
  1369 => x"81b72d85",
  1370 => x"1480f52d",
  1371 => x"73708105",
  1372 => x"5581b72d",
  1373 => x"871480f5",
  1374 => x"2d737081",
  1375 => x"055581b7",
  1376 => x"2d891480",
  1377 => x"f52d7370",
  1378 => x"81055581",
  1379 => x"b72d8e14",
  1380 => x"80f52d73",
  1381 => x"70810555",
  1382 => x"81b72d90",
  1383 => x"1480f52d",
  1384 => x"73708105",
  1385 => x"5581b72d",
  1386 => x"921480f5",
  1387 => x"2d737081",
  1388 => x"055581b7",
  1389 => x"2d941480",
  1390 => x"f52d7370",
  1391 => x"81055581",
  1392 => x"b72d9614",
  1393 => x"80f52d73",
  1394 => x"70810555",
  1395 => x"81b72d98",
  1396 => x"1480f52d",
  1397 => x"73708105",
  1398 => x"5581b72d",
  1399 => x"9c1480f5",
  1400 => x"2d737081",
  1401 => x"055581b7",
  1402 => x"2d9e1480",
  1403 => x"f52d7381",
  1404 => x"b72d77b9",
  1405 => x"9c0c8053",
  1406 => x"72bad80c",
  1407 => x"02a0050d",
  1408 => x"0402cc05",
  1409 => x"0d7e605e",
  1410 => x"5a800b80",
  1411 => x"c1fc0880",
  1412 => x"c2800859",
  1413 => x"5c568058",
  1414 => x"80c1dc08",
  1415 => x"782e81b0",
  1416 => x"38778f06",
  1417 => x"a0175754",
  1418 => x"738f38bb",
  1419 => x"cc527651",
  1420 => x"811757a0",
  1421 => x"812dbbcc",
  1422 => x"56807680",
  1423 => x"f52d5654",
  1424 => x"74742e83",
  1425 => x"38815474",
  1426 => x"81e52e80",
  1427 => x"f7388170",
  1428 => x"7506555c",
  1429 => x"73802e80",
  1430 => x"eb388b16",
  1431 => x"80f52d98",
  1432 => x"06597880",
  1433 => x"df388b53",
  1434 => x"7c527551",
  1435 => x"a1a12dba",
  1436 => x"d80880d0",
  1437 => x"389c1608",
  1438 => x"51aee92d",
  1439 => x"bad80884",
  1440 => x"1b0c9a16",
  1441 => x"80e02d51",
  1442 => x"af992dba",
  1443 => x"d808bad8",
  1444 => x"08881c0c",
  1445 => x"bad80855",
  1446 => x"5580c1d8",
  1447 => x"08802e98",
  1448 => x"38941680",
  1449 => x"e02d51af",
  1450 => x"992dbad8",
  1451 => x"08902b83",
  1452 => x"fff00a06",
  1453 => x"70165154",
  1454 => x"73881b0c",
  1455 => x"787a0c7b",
  1456 => x"54ae8904",
  1457 => x"81185880",
  1458 => x"c1dc0878",
  1459 => x"26fed238",
  1460 => x"80c1d808",
  1461 => x"802eb038",
  1462 => x"7a51a8dd",
  1463 => x"2dbad808",
  1464 => x"bad80880",
  1465 => x"fffffff8",
  1466 => x"06555b73",
  1467 => x"80ffffff",
  1468 => x"f82e9438",
  1469 => x"bad808fe",
  1470 => x"0580c1d0",
  1471 => x"082980c1",
  1472 => x"e4080557",
  1473 => x"ac960480",
  1474 => x"5473bad8",
  1475 => x"0c02b405",
  1476 => x"0d0402f4",
  1477 => x"050d7470",
  1478 => x"08810571",
  1479 => x"0c700880",
  1480 => x"c1d40806",
  1481 => x"5353718e",
  1482 => x"38881308",
  1483 => x"51a8dd2d",
  1484 => x"bad80888",
  1485 => x"140c810b",
  1486 => x"bad80c02",
  1487 => x"8c050d04",
  1488 => x"02f0050d",
  1489 => x"75881108",
  1490 => x"fe0580c1",
  1491 => x"d0082980",
  1492 => x"c1e40811",
  1493 => x"720880c1",
  1494 => x"d4080605",
  1495 => x"79555354",
  1496 => x"54a0812d",
  1497 => x"0290050d",
  1498 => x"0402f405",
  1499 => x"0d747088",
  1500 => x"2a83fe80",
  1501 => x"06707298",
  1502 => x"2a077288",
  1503 => x"2b87fc80",
  1504 => x"80067398",
  1505 => x"2b81f00a",
  1506 => x"06717307",
  1507 => x"07bad80c",
  1508 => x"56515351",
  1509 => x"028c050d",
  1510 => x"0402f805",
  1511 => x"0d028e05",
  1512 => x"80f52d74",
  1513 => x"882b0770",
  1514 => x"83ffff06",
  1515 => x"bad80c51",
  1516 => x"0288050d",
  1517 => x"0402f405",
  1518 => x"0d747678",
  1519 => x"53545280",
  1520 => x"71259738",
  1521 => x"72708105",
  1522 => x"5480f52d",
  1523 => x"72708105",
  1524 => x"5481b72d",
  1525 => x"ff115170",
  1526 => x"eb388072",
  1527 => x"81b72d02",
  1528 => x"8c050d04",
  1529 => x"02e8050d",
  1530 => x"77568070",
  1531 => x"56547376",
  1532 => x"24b33880",
  1533 => x"c1dc0874",
  1534 => x"2eab3873",
  1535 => x"51a9ce2d",
  1536 => x"bad808ba",
  1537 => x"d8080981",
  1538 => x"0570bad8",
  1539 => x"08079f2a",
  1540 => x"77058117",
  1541 => x"57575353",
  1542 => x"74762489",
  1543 => x"3880c1dc",
  1544 => x"087426d7",
  1545 => x"3872bad8",
  1546 => x"0c029805",
  1547 => x"0d0402f0",
  1548 => x"050dbad4",
  1549 => x"081651af",
  1550 => x"e42dbad8",
  1551 => x"08802e9c",
  1552 => x"388b53ba",
  1553 => x"d80852bf",
  1554 => x"cc51afb5",
  1555 => x"2d80c288",
  1556 => x"08547380",
  1557 => x"2e8638bf",
  1558 => x"cc51732d",
  1559 => x"0290050d",
  1560 => x"0402dc05",
  1561 => x"0d80705a",
  1562 => x"5574bad4",
  1563 => x"0825b138",
  1564 => x"80c1dc08",
  1565 => x"752ea938",
  1566 => x"7851a9ce",
  1567 => x"2dbad808",
  1568 => x"09810570",
  1569 => x"bad80807",
  1570 => x"9f2a7605",
  1571 => x"811b5b56",
  1572 => x"5474bad4",
  1573 => x"08258938",
  1574 => x"80c1dc08",
  1575 => x"7926d938",
  1576 => x"80557880",
  1577 => x"c1dc0827",
  1578 => x"81d13878",
  1579 => x"51a9ce2d",
  1580 => x"bad80880",
  1581 => x"2e81a538",
  1582 => x"bad8088b",
  1583 => x"0580f52d",
  1584 => x"70842a70",
  1585 => x"81067710",
  1586 => x"78842bbf",
  1587 => x"cc0b80f5",
  1588 => x"2d5c5c53",
  1589 => x"51555673",
  1590 => x"802e80c8",
  1591 => x"38741682",
  1592 => x"2bb39f0b",
  1593 => x"b9a8120c",
  1594 => x"54777531",
  1595 => x"1080c28c",
  1596 => x"11555690",
  1597 => x"74708105",
  1598 => x"5681b72d",
  1599 => x"a07481b7",
  1600 => x"2d7681ff",
  1601 => x"06811658",
  1602 => x"5473802e",
  1603 => x"89389c53",
  1604 => x"bfcc52b2",
  1605 => x"9c048b53",
  1606 => x"bad80852",
  1607 => x"80c28e16",
  1608 => x"51b2d404",
  1609 => x"7416822b",
  1610 => x"b0ae0bb9",
  1611 => x"a8120c54",
  1612 => x"7681ff06",
  1613 => x"81165854",
  1614 => x"73802e89",
  1615 => x"389c53bf",
  1616 => x"cc52b2cb",
  1617 => x"048b53ba",
  1618 => x"d8085277",
  1619 => x"75311080",
  1620 => x"c28c0551",
  1621 => x"7655afb5",
  1622 => x"2db2f004",
  1623 => x"74902975",
  1624 => x"31701080",
  1625 => x"c28c0551",
  1626 => x"54bad808",
  1627 => x"7481b72d",
  1628 => x"81195974",
  1629 => x"8b24a338",
  1630 => x"b1a20474",
  1631 => x"90297531",
  1632 => x"701080c2",
  1633 => x"8c058c77",
  1634 => x"31575154",
  1635 => x"807481b7",
  1636 => x"2d9e14ff",
  1637 => x"16565474",
  1638 => x"f33802a4",
  1639 => x"050d0402",
  1640 => x"fc050dba",
  1641 => x"d4081351",
  1642 => x"afe42dba",
  1643 => x"d808802e",
  1644 => x"8838bad8",
  1645 => x"0851a1df",
  1646 => x"2d800bba",
  1647 => x"d40cb0e1",
  1648 => x"2d8ee72d",
  1649 => x"0284050d",
  1650 => x"0402fc05",
  1651 => x"0d725170",
  1652 => x"fd2ead38",
  1653 => x"70fd248a",
  1654 => x"3870fc2e",
  1655 => x"80c438b4",
  1656 => x"aa0470fe",
  1657 => x"2eb13870",
  1658 => x"ff2e0981",
  1659 => x"06bc38ba",
  1660 => x"d4085170",
  1661 => x"802eb338",
  1662 => x"ff11bad4",
  1663 => x"0cb4aa04",
  1664 => x"bad408f0",
  1665 => x"0570bad4",
  1666 => x"0c517080",
  1667 => x"259c3880",
  1668 => x"0bbad40c",
  1669 => x"b4aa04ba",
  1670 => x"d4088105",
  1671 => x"bad40cb4",
  1672 => x"aa04bad4",
  1673 => x"089005ba",
  1674 => x"d40cb0e1",
  1675 => x"2d8ee72d",
  1676 => x"0284050d",
  1677 => x"0402fc05",
  1678 => x"0d800bba",
  1679 => x"d40cb0e1",
  1680 => x"2d8ddf2d",
  1681 => x"bad808ba",
  1682 => x"c40cb9a0",
  1683 => x"5190822d",
  1684 => x"0284050d",
  1685 => x"047180c2",
  1686 => x"880c0400",
  1687 => x"00ffffff",
  1688 => x"ff00ffff",
  1689 => x"ffff00ff",
  1690 => x"ffffff00",
  1691 => x"52657365",
  1692 => x"74204e45",
  1693 => x"53000000",
  1694 => x"5363616e",
  1695 => x"6c696e65",
  1696 => x"73000000",
  1697 => x"48513258",
  1698 => x"2046696c",
  1699 => x"74657200",
  1700 => x"33206f72",
  1701 => x"20362062",
  1702 => x"7574746f",
  1703 => x"6e206a6f",
  1704 => x"79737469",
  1705 => x"636b0000",
  1706 => x"50312053",
  1707 => x"656c6563",
  1708 => x"74000000",
  1709 => x"50312053",
  1710 => x"74617274",
  1711 => x"00000000",
  1712 => x"4c6f6164",
  1713 => x"20524f4d",
  1714 => x"20100000",
  1715 => x"45786974",
  1716 => x"00000000",
  1717 => x"524f4d20",
  1718 => x"6c6f6164",
  1719 => x"696e6720",
  1720 => x"6661696c",
  1721 => x"65640000",
  1722 => x"4f4b0000",
  1723 => x"496e6974",
  1724 => x"69616c69",
  1725 => x"7a696e67",
  1726 => x"20534420",
  1727 => x"63617264",
  1728 => x"0a000000",
  1729 => x"16200000",
  1730 => x"14200000",
  1731 => x"15200000",
  1732 => x"53442069",
  1733 => x"6e69742e",
  1734 => x"2e2e0a00",
  1735 => x"53442063",
  1736 => x"61726420",
  1737 => x"72657365",
  1738 => x"74206661",
  1739 => x"696c6564",
  1740 => x"210a0000",
  1741 => x"53444843",
  1742 => x"20657272",
  1743 => x"6f72210a",
  1744 => x"00000000",
  1745 => x"57726974",
  1746 => x"65206661",
  1747 => x"696c6564",
  1748 => x"0a000000",
  1749 => x"52656164",
  1750 => x"20666169",
  1751 => x"6c65640a",
  1752 => x"00000000",
  1753 => x"43617264",
  1754 => x"20696e69",
  1755 => x"74206661",
  1756 => x"696c6564",
  1757 => x"0a000000",
  1758 => x"46415431",
  1759 => x"36202020",
  1760 => x"00000000",
  1761 => x"46415433",
  1762 => x"32202020",
  1763 => x"00000000",
  1764 => x"4e6f2070",
  1765 => x"61727469",
  1766 => x"74696f6e",
  1767 => x"20736967",
  1768 => x"0a000000",
  1769 => x"42616420",
  1770 => x"70617274",
  1771 => x"0a000000",
  1772 => x"4261636b",
  1773 => x"00000000",
  1774 => x"00000002",
  1775 => x"00000002",
  1776 => x"00001a6c",
  1777 => x"0000034e",
  1778 => x"00000001",
  1779 => x"00001a78",
  1780 => x"00000000",
  1781 => x"00000001",
  1782 => x"00001a84",
  1783 => x"00000001",
  1784 => x"00000001",
  1785 => x"00001a90",
  1786 => x"00000002",
  1787 => x"00000002",
  1788 => x"00001aa8",
  1789 => x"00000362",
  1790 => x"00000002",
  1791 => x"00001ab4",
  1792 => x"00000376",
  1793 => x"00000002",
  1794 => x"00001ac0",
  1795 => x"00001a35",
  1796 => x"00000002",
  1797 => x"00001acc",
  1798 => x"000006f9",
  1799 => x"00000000",
  1800 => x"00000000",
  1801 => x"00000000",
  1802 => x"00000004",
  1803 => x"00001ad4",
  1804 => x"00001c28",
  1805 => x"00000004",
  1806 => x"00001ae8",
  1807 => x"00001bbc",
  1808 => x"00000000",
  1809 => x"00000000",
  1810 => x"00000000",
  1811 => x"00000000",
  1812 => x"00000000",
  1813 => x"00000000",
  1814 => x"00000000",
  1815 => x"00000000",
  1816 => x"00000000",
  1817 => x"00000000",
  1818 => x"00000000",
  1819 => x"00000000",
  1820 => x"00000000",
  1821 => x"00000000",
  1822 => x"00000000",
  1823 => x"00000000",
  1824 => x"00000000",
  1825 => x"00000000",
  1826 => x"00000000",
  1827 => x"00000000",
  1828 => x"00000000",
  1829 => x"00000000",
  1830 => x"00000000",
  1831 => x"00000000",
  1832 => x"00000002",
  1833 => x"0000210c",
  1834 => x"0000182e",
  1835 => x"00000002",
  1836 => x"0000212a",
  1837 => x"0000182e",
  1838 => x"00000002",
  1839 => x"00002148",
  1840 => x"0000182e",
  1841 => x"00000002",
  1842 => x"00002166",
  1843 => x"0000182e",
  1844 => x"00000002",
  1845 => x"00002184",
  1846 => x"0000182e",
  1847 => x"00000002",
  1848 => x"000021a2",
  1849 => x"0000182e",
  1850 => x"00000002",
  1851 => x"000021c0",
  1852 => x"0000182e",
  1853 => x"00000002",
  1854 => x"000021de",
  1855 => x"0000182e",
  1856 => x"00000002",
  1857 => x"000021fc",
  1858 => x"0000182e",
  1859 => x"00000002",
  1860 => x"0000221a",
  1861 => x"0000182e",
  1862 => x"00000002",
  1863 => x"00002238",
  1864 => x"0000182e",
  1865 => x"00000002",
  1866 => x"00002256",
  1867 => x"0000182e",
  1868 => x"00000002",
  1869 => x"00002274",
  1870 => x"0000182e",
  1871 => x"00000004",
  1872 => x"00001bb0",
  1873 => x"00000000",
  1874 => x"00000000",
  1875 => x"00000000",
  1876 => x"000019c9",
  1877 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;

